library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.ALL;

package geometryPackage is

type romArray is array (0 to 132-1) of integer;
type incArray is array (0 to 2) of integer;

-- All the notes periods in integers where mod4 == 0
constant T : romArray := (12231220, 11544732, 10896776, 10285188, 9707924, 9163060, 8648780, 8163360, 7705184, 7272728, 6864540, 6479264, 6115608, 5772368, 5448388, 5142592, 4853964, 4581532, 4324388, 4081680, 3852592, 3636364, 3432268, 3239632, 3057804, 2886184, 2724192, 2571296, 2426980, 2290764, 2162192, 2040840, 1926296, 1818180, 1716136, 1619816, 1528900, 1443092, 1362096, 1285648, 1213488, 1145380, 1081096, 1020420, 963148, 909088, 858068, 809908, 764452, 721544, 681048, 642824, 606744, 572692, 540548, 510208, 481572, 454544, 429032, 404952, 382224, 360772, 340524, 321412, 303372, 286344, 270272, 255104, 240788, 227272, 214516, 202476, 191112, 180384, 170260, 160704, 151684, 143172, 135136, 127552, 120392, 113636, 107256, 101236, 95556, 90192, 85132, 80352, 75844, 71584, 67568, 63776, 60196, 56816, 53628, 50620, 47776, 45096, 42564, 40176, 37920, 35792, 33784, 31888, 30096, 28408, 26812, 25308, 23888, 22548, 21280, 20088, 18960, 17896, 16892, 15944, 15048, 14204, 13408, 12652, 11944, 11272, 10640, 10044, 9480, 8948, 8444, 7972, 7524, 7100, 6704, 6328);
-- All the periods for their respective sampling frequencies
--constant F_s : romArray := (611561, 577237, 544839, 514259, 485396, 458153, 432439, 408168, 385259, 363636, 343227, 323963, 305781, 288618, 272419, 257130, 242698, 229077, 216219, 204084, 192630, 181818, 171614, 161982, 152890, 144309, 136210, 128565, 121349, 114538, 108110, 102042, 96315, 90909, 85807, 80991, 76445, 72155, 68105, 64282, 60675, 57269, 54055, 51021, 48157, 45455, 42903, 40495, 38223, 36077, 34052, 32141, 30337, 28635, 27027, 25511, 24079, 22727, 21452, 20248, 19111, 18039, 17026, 16071, 15169, 14317, 13514, 12755, 12039, 11364, 10726, 10124, 9556, 9019, 8513, 8035, 7584, 7159, 6757, 6378, 6020, 5682, 5363, 5062, 4778, 4510, 4257, 4018, 3792, 3579, 3378, 3189, 3010, 2841, 2681, 2531, 2389, 2255, 2128, 2009, 1896, 1790, 1689, 1594, 1505, 1420, 1341, 1265, 1194, 1127, 1064, 1004, 948, 895, 845, 797, 752, 710, 670, 633, 597, 564, 532, 502, 474, 447, 422, 399, 376, 355, 335, 316);
constant F_s : romArray := (407707, 384824, 363226, 342840, 323598, 305435, 288293, 272112, 256840, 242424, 228818, 215975, 203854, 192412, 181613, 171420, 161799, 152718, 144146, 136056, 128420, 121212, 114409, 107988, 101927, 96206, 90806, 85710, 80899, 76359, 72073, 68028, 64210, 60606, 57205, 53994, 50963, 48103, 45403, 42855, 40450, 38179, 36037, 34014, 32105, 30303, 28602, 26997, 25482, 24052, 22702, 21427, 20225, 19090, 18018, 17007, 16052, 15152, 14301, 13498, 12741, 12026, 11351, 10714, 10112, 9545, 9009, 8504, 8026, 7576, 7151, 6749, 6370, 6013, 5675, 5357, 5056, 4772, 4505, 4252, 4013, 3788, 3575, 3375, 3185, 3006, 2838, 2678, 2528, 2386, 2252, 2126, 2007, 1894, 1788, 1687, 1593, 1503, 1419, 1339, 1264, 1193, 1126, 1063, 1003, 947, 894, 844, 796, 752, 709, 670, 632, 597, 563, 531, 502, 473, 447, 422, 398, 376, 355, 335, 316, 298, 282, 266, 251, 237, 223, 211);
-- The incrementation at every sampling point
constant inc : incArray := (18078, 9039, 16383);

-- Declare functions
function getT (input : integer) return integer;
function getFs (input : integer) return integer;
function getInc (input : integer) return integer;

end geometryPackage;

package body geometryPackage is

    function getT (input : integer) return integer is
    begin
        return T(input);
    end getT;
    
    function getFs (input : integer) return integer is
    begin
        return F_s(input);
    end getFs;
    
    function getInc (input : integer) return integer is
    begin
        return inc(input);
    end getInc;

end geometryPackage;
