library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.ALL;

package geometryPackage is

type romArray is array (0 to 132-1) of integer;

-- All the notes periods in integers where mod4 == 0
constant T : romArray := (12231220, 11544732, 10896776, 10285188, 9707924, 9163060, 8648780, 8163360, 7705184, 7272728, 6864540, 6479264, 6115608, 5772368, 5448388, 5142592, 4853964, 4581532, 4324388, 4081680, 3852592, 3636364, 3432268, 3239632, 3057804, 2886184, 2724192, 2571296, 2426980, 2290764, 2162192, 2040840, 1926296, 1818180, 1716136, 1619816, 1528900, 1443092, 1362096, 1285648, 1213488, 1145380, 1081096, 1020420, 963148, 909088, 858068, 809908, 764452, 721544, 681048, 642824, 606744, 572692, 540548, 510208, 481572, 454544, 429032, 404952, 382224, 360772, 340524, 321412, 303372, 286344, 270272, 255104, 240788, 227272, 214516, 202476, 191112, 180384, 170260, 160704, 151684, 143172, 135136, 127552, 120392, 113636, 107256, 101236, 95556, 90192, 85132, 80352, 75844, 71584, 67568, 63776, 60196, 56816, 53628, 50620, 47776, 45096, 42564, 40176, 37920, 35792, 33784, 31888, 30096, 28408, 26812, 25308, 23888, 22548, 21280, 20088, 18960, 17896, 16892, 15944, 15048, 14204, 13408, 12652, 11944, 11272, 10640, 10044, 9480, 8948, 8444, 7972, 7524, 7100, 6704, 6328);
-- All the periods for their respective sampling frequencies
constant F_s : romArray := (1223122, 1154473, 1089678, 1028519, 970793, 916306, 864878, 816336, 770519, 727273, 686454, 647926, 611561, 577237, 544839, 514259, 485396, 458153, 432439, 408168, 385259, 363636, 343227, 323963, 305781, 288618, 272419, 257130, 242698, 229077, 216219, 204084, 192630, 181818, 171614, 161982, 152890, 144309, 136210, 128565, 121349, 114538, 108110, 102042, 96315, 90909, 85807, 80991, 76445, 72155, 68105, 64282, 60675, 57269, 54055, 51021, 48157, 45455, 42903, 40495, 38223, 36077, 34052, 32141, 30337, 28635, 27027, 25511, 24079, 22727, 21452, 20248, 19111, 18039, 17026, 16071, 15169, 14317, 13514, 12755, 12039, 11364, 10726, 10124, 9556, 9019, 8513, 8035, 7584, 7159, 6757, 6378, 6020, 5682, 5363, 5062, 4778, 4510, 4257, 4018, 3792, 3579, 3378, 3189, 3010, 2841, 2681, 2531, 2389, 2255, 2128, 2009, 1896, 1790, 1689, 1594, 1505, 1420, 1341, 1265, 1194, 1127, 1064, 1004, 948, 895, 845, 797, 752, 710, 670, 633);
-- The incrementation at every sampling point
constant inc : romArray := (3, 3, 3, 4, 4, 4, 4, 5, 5, 5, 6, 6, 6, 7, 7, 8, 8, 9, 9, 10, 10, 11, 12, 12, 13, 14, 15, 16, 17, 18, 19, 20, 21, 23, 24, 25, 27, 29, 30, 32, 34, 36, 38, 41, 43, 46, 48, 51, 54, 58, 61, 65, 69, 73, 77, 82, 87, 92, 97, 103, 109, 116, 123, 130, 138, 146, 155, 164, 174, 184, 195, 207, 219, 232, 246, 260, 276, 292, 310, 328, 348, 369, 391, 414, 438, 465, 492, 522, 553, 585, 620, 657, 696, 738, 782, 828, 877, 930, 985, 1043, 1106, 1171, 1241, 1315, 1393, 1476, 1564, 1657, 1755, 1860, 1971, 2087, 2212, 2343, 2483, 2631, 2786, 2953, 3127, 3315, 3512, 3721, 3942, 4177, 4424, 4686, 4963, 5262, 5577, 5907, 6260, 6626);

-- Declare functions
function getT (input : integer) return integer;
function getFs (input : integer) return integer;
function getInc (input : integer) return integer;

end geometryPackage;

package body geometryPackage is

    function getT (input : integer) return integer is
    begin
        return T(input);
    end getT;
    
    function getFs (input : integer) return integer is
    begin
        return F_s(input);
    end getFs;
    
    function getInc (input : integer) return integer is
    begin
        return inc(input);
    end getInc;

end geometryPackage;
