library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity sine is
end sine;

architecture Behavioral of sine is

begin


end Behavioral;

